--Commit 3 by Bren