--Commit 4 by Brent