--Commit 3 by Brent